`define TYPE_I 7'b0010011